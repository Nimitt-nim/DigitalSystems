module Decoder(
    input [4:0]A;
    output [31:0]OUT;
);

always @(*)
    OUT[0] = (~A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4]);
    OUT[1] = (A[0] & ~A[1] & ~A[2] & ~A[3] & ~A[4]);
    OUT[2] = (~A[0] & A[1] & ~A[2] & ~A[3] & ~A[4]);
    OUT[3] = (A[0] & A[1] & ~A[2] & ~A[3] & ~A[4]);
    OUT[4] = (~A[0] & ~A[1] & A[2] & ~A[3] & ~A[4]);
    OUT[5] = (A[0] & ~A[1] & A[2] & ~A[3] & ~A[4]);
    OUT[6] = (~A[0] & A[1] & A[2] & ~A[3] & ~A[4]);
    OUT[7] = (A[0] & A[1] & A[2] & ~A[3] & ~A[4]);
    OUT[8] = (~A[0] & ~A[1] & ~A[2] & A[3] & ~A[4]);
    OUT[9] = (A[0] & ~A[1] & ~A[2] & A[3] & ~A[4]);
    OUT[10] = (~A[0] & A[1] & ~A[2] & A[3] & ~A[4]);
    OUT[11] = (A[0] & A[1] & ~A[2] & A[3] & ~A[4]);
    OUT[12] = (~A[0] & ~A[1] & A[2] & A[3] & ~A[4]);
    OUT[13] = (A[0] & ~A[1] & A[2] & A[3] & ~A[4]);
    OUT[14] = (~A[0] & A[1] & A[2] & A[3] & ~A[4]);
    OUT[15] = (A[0] & A[1] & A[2] & A[3] & ~A[4]);

    OUT[16] = (~A[0] & ~A[1] & ~A[2] & ~A[3] & A[4]);
    OUT[17] = (A[0] & ~A[1] & ~A[2] & ~A[3] & A[4]);
    OUT[18] = (~A[0] & A[1] & ~A[2] & ~A[3] & A[4]);
    OUT[19] = (A[0] & A[1] & ~A[2] & ~A[3] & A[4]);
    OUT[20] = (~A[0] & ~A[1] & A[2] & ~A[3] & A[4]);
    OUT[21] = (A[0] & ~A[1] & A[2] & ~A[3] & A[4]);
    OUT[22] = (~A[0] & A[1] & A[2] & ~A[3] & A[4]);
    OUT[23] = (A[0] & A[1] & A[2] & ~A[3] & A[4]);
    OUT[24] = (~A[0] & ~A[1] & ~A[2] & A[3] & A[4]);
    OUT[25] = (A[0] & ~A[1] & ~A[2] & A[3] & A[4]);
    OUT[26] = (~A[0] & A[1] & ~A[2] & A[3] & A[4]);
    OUT[27] = (A[0] & A[1] & ~A[2] & A[3] & A[4]);
    OUT[28] = (~A[0] & ~A[1] & A[2] & A[3] & A[4]);
    OUT[29] = (A[0] & ~A[1] & A[2] & A[3] & A[4]);
    OUT[30] = (~A[0] & A[1] & A[2] & A[3] & A[4]);
    OUT[31] = (A[0] & A[1] & A[2] & A[3] & A[4]);

    
endmodule