module Decoder(
    input [4:0]R;
    output [31:0]OUT3;
);

always @(*)
    OUT3[0] = (R[0] || R[1] || R[2] || R[3] || R[4]);
    OUT3[1] = (R[0] || R[1] || R[2] || R[3] || R[4]);
    OUT3[2] = (R[1] || R[2] || R[3] || R[4]);
    OUT3[3] = ((R[0] & R[1]) || R[2] || R[3] || R[4]);
    OUT3[4] = (R[1] || R[2] || R[3] || R[4]);
    OUT3[5] = ((R[0] & R[2]) || R[3] || R[4]);
    OUT3[6] = ((R[1] & R[2]) || R[2] || R[3] || R[4]);
    OUT3[7] = ((R[0] & R[1] & R[2]) || R[2] || R[3] || R[4]);
    OUT3[8] = (R[3] || R[4]);
    OUT3[9] = (R[0] & ~R[1] & ~R[2] & R[3] & ~R[4]);
    OUT3[10] = (~R[0] & R[1] & ~R[2] & R[3] & ~R[4]);
    OUT3[11] = (R[0] & R[1] & ~R[2] & R[3] & ~R[4]);
    OUT3[12] = (~R[0] & ~R[1] & R[2] & R[3] & ~R[4]);
    OUT3[13] = (R[0] & ~R[1] & R[2] & R[3] & ~R[4]);
    OUT3[14] = (~R[0] & R[1] & R[2] & R[3] & ~R[4]);
    OUT3[15] = (R[0] & R[1] & R[2] & R[3] & ~R[4]);

    OUT3[16] = (R[4]);
    OUT3[17] = (R[4] & ( R[0] || R[1] || R[2] || R[3]));
    OUT3[18] = (R[4] & ( R[0] || R[1] || R[2] || R[3]))
    OUT3[19] = (R[0] & R[1] & ~R[2] & ~R[3] & R[4]);
    OUT3[20] = (~R[0] & ~R[1] & R[2] & ~R[3] & R[4]);
    OUT3[21] = (R[0] & ~R[1] & R[2] & ~R[3] & R[4]);
    OUT3[22] = (~R[0] & R[1] & R[2] & ~R[3] & R[4]);
    OUT3[23] = (R[0] & R[1] & R[2] & ~R[3] & R[4]);
    OUT3[24] = (~R[0] & ~R[1] & ~R[2] & R[3] & R[4]);
    OUT3[25] = (R[0] & ~R[1] & ~R[2] & R[3] & R[4]);
    OUT3[26] = (~R[0] & R[1] & ~R[2] & R[3] & R[4]);
    OUT3[27] = (R[0] & R[1] & ~R[2] & R[3] & R[4]);
    OUT3[28] = (~R[0] & ~R[1] & R[2] & R[3] & R[4]);
    OUT3[29] = (R[0] & ~R[1] & R[2] & R[3] & R[4]);
    OUT3[30] = (OUT3[31]|| R[]);
    OUT3[31] = (~R[0] & ~R[1] & ~R[2] & ~R[3] & ~R[4]);

    
endmodule