module SmartMathTutor(
    input[4:0]R;
    input[9:2]S;
    output [31:0]OUT;
);

always @(*)
    begin
    // Decoder
    Rd[0] = (~R[0] & ~R[1] & ~R[2] & ~R[3] & ~R[4]);
    Rd[1] = (R[0] & ~R[1] & ~R[2] & ~R[3] & ~R[4]);
    Rd[2] = (~R[0] & R[1] & ~R[2] & ~R[3] & ~R[4]);
    Rd[3] = (R[0] & R[1] & ~R[2] & ~R[3] & ~R[4]);
    Rd[4] = (~R[0] & ~R[1] & R[2] & ~R[3] & ~R[4]);
    Rd[5] = (R[0] & ~R[1] & R[2] & ~R[3] & ~R[4]);
    Rd[6] = (~R[0] & R[1] & R[2] & ~R[3] & ~R[4]);
    Rd[7] = (R[0] & R[1] & R[2] & ~R[3] & ~R[4]);
    Rd[8] = (~R[0] & ~R[1] & ~R[2] & R[3] & ~R[4]);
    Rd[9] = (R[0] & ~R[1] & ~R[2] & R[3] & ~R[4]);
    Rd[10] = (~R[0] & R[1] & ~R[2] & R[3] & ~R[4]);
    Rd[11] = (R[0] & R[1] & ~R[2] & R[3] & ~R[4]);
    Rd[12] = (~R[0] & ~R[1] & R[2] & R[3] & ~R[4]);
    Rd[13] = (R[0] & ~R[1] & R[2] & R[3] & ~R[4]);
    Rd[14] = (~R[0] & R[1] & R[2] & R[3] & ~R[4]);
    Rd[15] = (R[0] & R[1] & R[2] & R[3] & ~R[4]);
    Rd[16] = (~R[0] & ~R[1] & ~R[2] & ~R[3] & R[4]);
    Rd[17] = (R[0] & ~R[1] & ~R[2] & ~R[3] & R[4]);
    Rd[18] = (~R[0] & R[1] & ~R[2] & ~R[3] & R[4]);
    Rd[19] = (R[0] & R[1] & ~R[2] & ~R[3] & R[4]);
    Rd[20] = (~R[0] & ~R[1] & R[2] & ~R[3] & R[4]);
    Rd[21] = (R[0] & ~R[1] & R[2] & ~R[3] & R[4]);
    Rd[22] = (~R[0] & R[1] & R[2] & ~R[3] & R[4]);
    Rd[23] = (R[0] & R[1] & R[2] & ~R[3] & R[4]);
    Rd[24] = (~R[0] & ~R[1] & ~R[2] & R[3] & R[4]);
    Rd[25] = (R[0] & ~R[1] & ~R[2] & R[3] & R[4]);
    Rd[26] = (~R[0] & R[1] & ~R[2] & R[3] & R[4]);
    Rd[27] = (R[0] & R[1] & ~R[2] & R[3] & R[4]);
    Rd[28] = (~R[0] & ~R[1] & R[2] & R[3] & R[4]);
    Rd[29] = (R[0] & ~R[1] & R[2] & R[3] & R[4]);
    Rd[30] = (~R[0] & R[1] & R[2] & R[3] & R[4]);
    Rd[31] = (R[0] & R[1] & R[2] & R[3] & R[4]);

    // Range
    Rc[31] = (~R[0] & ~R[1] & ~R[2] & ~R[3] & ~R[4]);
    Rc[30] = (Rc[31] | Rd[30]);
    Rc[29] = (Rc[30] | Rd[29]);
    Rc[28] = (Rc[29] | Rd[28]);
    Rc[27] = (Rc[28] | Rd[27]);
    Rc[26] = (Rc[27] | Rd[26]);
    Rc[25] = (Rc[26] | Rd[25]);
    Rc[24] = (Rc[25] | Rd[24]);
    Rc[23] = (Rc[24] | Rd[23]);
    Rc[22] = (Rc[23] | Rd[22]);
    Rc[21] = (Rc[22] | Rd[21]);
    Rc[20] = (Rc[21] | Rd[20]);
    Rc[19] = (Rc[20] | Rd[19]);
    Rc[18] = (Rc[19] | Rd[18]);
    Rc[17] = (Rc[18] | Rd[17]);
    Rc[16] = (Rc[17] | Rd[16]);
    Rc[15] = (Rc[16] | Rd[15]);
    Rc[14] = (Rc[15] | Rd[14]);
    Rc[13] = (Rc[14] | Rd[13]);
    Rc[12] = (Rc[13] | Rd[12]);
    Rc[11] = (Rc[12] | Rd[11]);
    Rc[10] = (Rc[11] | Rd[10]);
    Rc[9] = (Rc[10]  | Rd[9]);
    Rc[8] = (Rc[9] | Rd[8]);
    Rc[7] = (Rc[8] | Rd[7]);
    Rc[6] = (Rc[7] | Rd[6]);
    Rc[5] = (Rc[6] | Rd[5]);
    Rc[4] = (Rc[5] | Rd[4]);
    Rc[3] = (Rc[4] | Rd[3]);
    Rc[2] = (Rc[3] | Rd[2]);
    Rc[1] = (Rc[2] | Rd[1]);
    Rc[0] = (Rc[1] | Rd[0]);


    // creating the final out put array
    OUT[0] =   1;
    OUT[1] =   0;
    OUT[2] =   S[2] &&  Rc[2];
    OUT[3] =   S[3] &&  Rc[3];
    OUT[4] =   S[2] | S[4] &&  Rc[4];
    OUT[5] =   S[5] &&  Rc[5];
    OUT[6] =   S[2] | S[3] &&  Rc[6];
    OUT[7] =   S[7] &&  Rc[7];
    OUT[8] =   S[2] | S[4] | S[8] &&  Rc[8];
    OUT[9] =   S[3] | S[9] &&  Rc[9];
    OUT[10] =  S[2] | S[5] &&  Rc[10];
    OUT[11] =  0;
    OUT[12] =  S[2] | S[3] | S[4] | S[6]  &&  Rc[12];
    OUT[13] =  0;
    OUT[14] =  S[2] | S[7] &&  Rc[14];
    OUT[15] =  S[3] | S[5] &&  Rc[15];
    OUT[16] =  S[2] | S[4] | S[8] &&  Rc[16];
    OUT[17] =  0;
    OUT[18] =  S[2] | S[3] | S[6] | S[9] &&  Rc[18];
    OUT[19] =  0;
    OUT[20] =  S[2] | S[4] | S[5] &&  Rc[20];
    OUT[21] =  S[3] | S[7] | S[5] &&  Rc[21];
    OUT[22] =  S[2] &&  Rc[22];
    OUT[23] =  0;
    OUT[24] =  S[3] | S[7] | S[5] &&  Rc[24];
    OUT[25] =  S[5] &&  Rc[25];
    OUT[26] =  0;
    OUT[27] =  S[3] | S[9] &&  Rc[27];
    OUT[28] =  S[2] | S[4] | S[7] &&  Rc[28];
    OUT[29] =  0;
    OUT[30] =  S[2] | |S[3] | S[5] &&  Rc[30];
    OUT[31] =  0;
    end

endmodule